`timescale 1ns/100ps

module pipeline2(CLK, RESET, BRANCH, REG_DEST,MEM_TO_REG,ALU_SOURCE,MEM_READ,MEM_WRITE,IMMI_SEL, ALU_OP, OUT1, OUT2, PC_INCREMENT4,SIGN_EXTENDED, RD1, RD2, BUSY_WAIT,
BRANCH_OUT,REG_DEST_OUT,MEM_TO_REG_OUT,ALU_SOURCE_OUT,MEM_READ_OUT,MEM_WRITE_OUT,IMMI_SEL_OUT,ALU_OP_OUT,OUT1_OUT, OUT2_OUT, PC_INCREMENT4_OUT, SIGN_EXTENDED_OUT, RD1_OUT, RD2_OUT);
	input CLK, RESET, BRANCH,REG_DEST, REG_WRITE, BUSY_WAIT;
	input [1:0] MEM_TO_REG,ALU_SOURCE;
	input [2:0] MEM_READ,MEM_WRITE,IMMI_SEL;
	input [4:0] ALU_OP,RD1, RD2;
	input [31:0] OUT1, OUT2, PC_INCREMENT4, SIGN_EXTENDED;
	
	output reg BRANCH_OUT,REG_DEST_OUT, REG_WRITE_OUT;
	output reg [1:0] MEM_TO_REG_OUT,ALU_SOURCE_OUT;
	output reg [2:0] MEM_READ_OUT,MEM_WRITE_OUT,IMMI_SEL_OUT;
	output reg [4:0] ALU_OP_OUT,RD1_OUT,RD2_OUT;
	output reg [31:0] OUT1_OUT, OUT2_OUT, PC_INCREMENT4_OUT, SIGN_EXTENDED_OUT;
	
	always @(posedge CLK) begin
		if(!BUSY_WAIT) begin
			BRANCH_OUT = BRANCH;
			REG_DEST_OUT = REG_DEST;
			MEM_TO_REG_OUT = MEM_TO_REG;
			ALU_SOURCE_OUT = ALU_SOURCE;
			MEM_READ_OUT = MEM_READ;
			MEM_WRITE_OUT = MEM_WRITE;
			IMMI_SEL_OUT = IMMI_SEL;
			ALU_OP_OUT = ALU_OP;
			OUT1_OUT = OUT1;
			OUT2_OUT = OUT2;
			PC_INCREMENT4_OUT = PC_INCREMENT4;
			SIGN_EXTENDED_OUT = SIGN_EXTENDED;
			REG_WRITE_OUT = REG_WRITE;
		
		end
	end
endmodule